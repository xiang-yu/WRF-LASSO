netcdf force_template {
dimensions:
	Time = UNLIMITED ; // (0 currently)
	DateStrLen = 19 ;
	force_layers = 4;
variables:
	char Times(Time, DateStrLen) ;
	float Z_LS(Time, force_layers) ;
		Z_LS:FieldType = 104 ;
		Z_LS:MemoryOrder = "Z  " ;
		Z_LS:description = "height of forcing time series" ;
		Z_LS:units = "" ;
		Z_LS:stagger = "" ;
		Z_LS:_FillValue = -999.f ;
        float U_LS(Time, force_layers) ;
                U_LS:FieldType = 104 ;
                U_LS:MemoryOrder = "Z  " ;
                U_LS:description = "large scale zonal wind velocity" ;
                U_LS:units = "" ;
                U_LS:stagger = "" ;
                U_LS:_FillValue = -999.f ;
        float V_LS(Time, force_layers) ;
                V_LS:FieldType = 104 ;
                V_LS:MemoryOrder = "Z  " ;
                V_LS:description = "large scale meridional wind velocity" ;
                V_LS:units = "" ;
                V_LS:stagger = "" ;
                V_LS:_FillValue = -999.f ;
	float W_LS(Time, force_layers) ;
		W_LS:FieldType = 104 ;
		W_LS:MemoryOrder = "Z  " ;
		W_LS:description = "height of forcing time series" ;
		W_LS:units = "" ;
		W_LS:stagger = "" ;
		W_LS:_FillValue = -999.f ;
	float TH_ADV(Time, force_layers) ;
		TH_ADV:FieldType = 104 ;
		TH_ADV:MemoryOrder = "Z  " ;
		TH_ADV:description = "tendency of thermal adv" ;
		TH_ADV:units = "" ;
		TH_ADV:stagger = "" ;
		TH_ADV:_FillValue = -999.f ;
	float TH_RLX(Time, force_layers) ;
		TH_RLX:FieldType = 104 ;
		TH_RLX:MemoryOrder = "Z  " ;
		TH_RLX:description = "relaxation" ;
		TH_RLX:units = "" ;
		TH_RLX:stagger = "" ;
		TH_RLX:_FillValue = -999.f ;
	float QV_ADV(Time, force_layers) ;
		QV_ADV:FieldType = 104 ;
		QV_ADV:MemoryOrder = "Z  " ;
		QV_ADV:description = "tendency of qv adv" ;
		QV_ADV:units = "" ;
		QV_ADV:stagger = "" ;
		QV_ADV:_FillValue = -999.f ;
	float QV_RLX(Time, force_layers) ;
		QV_RLX:FieldType = 104 ;
		QV_RLX:MemoryOrder = "Z  " ;
		QV_RLX:description = "qv relaxation" ;
		QV_RLX:units = "" ;
		QV_RLX:stagger = "" ;
		QV_RLX:_FillValue = -999.f ;
	float Z_LS_TEND(Time, force_layers) ;
		Z_LS_TEND:FieldType = 104 ;
		Z_LS_TEND:MemoryOrder = "Z  " ;
		Z_LS_TEND:description = "height of forcing time series" ;
		Z_LS_TEND:units = "" ;
		Z_LS_TEND:stagger = "" ;
		Z_LS_TEND:_FillValue = -999.f ;
        float U_LS_TEND(Time, force_layers) ;
                U_LS_TEND:FieldType = 104 ;
                U_LS_TEND:MemoryOrder = "Z  " ;
                U_LS_TEND:description = "tendency of zonal wind" ;
                U_LS_TEND:units = "" ;
                U_LS_TEND:stagger = "" ;
                U_LS_TEND:_FillValue = -999.f ;
        float V_LS_TEND(Time, force_layers) ;
                V_LS_TEND:FieldType = 104 ;
                V_LS_TEND:MemoryOrder = "Z  " ;
                V_LS_TEND:description = "tendency of meridional wind" ;
                V_LS_TEND:units = "" ;
                V_LS_TEND:stagger = "" ;
                V_LS_TEND:_FillValue = -999.f ;
	float W_LS_TEND(Time, force_layers) ;
		W_LS_TEND:FieldType = 104 ;
		W_LS_TEND:MemoryOrder = "Z  " ;
		W_LS_TEND:description = "height of forcing time series" ;
		W_LS_TEND:units = "" ;
		W_LS_TEND:stagger = "" ;
		W_LS_TEND:_FillValue = -999.f ;
	float TH_ADV_TEND(Time, force_layers) ;
		TH_ADV_TEND:FieldType = 104 ;
		TH_ADV_TEND:MemoryOrder = "Z  " ;
		TH_ADV_TEND:description = "tendency of thermal adv" ;
		TH_ADV_TEND:units = "" ;
		TH_ADV_TEND:stagger = "" ;
		TH_ADV_TEND:_FillValue = -999.f ;
	float TH_RLX_TEND(Time, force_layers) ;
		TH_RLX_TEND:FieldType = 104 ;
		TH_RLX_TEND:MemoryOrder = "Z  " ;
		TH_RLX_TEND:description = "relaxation" ;
		TH_RLX_TEND:units = "" ;
		TH_RLX_TEND:stagger = "" ;
		TH_RLX_TEND:_FillValue = -999.f ;
	float QV_ADV_TEND(Time, force_layers) ;
		QV_ADV_TEND:FieldType = 104 ;
		QV_ADV_TEND:MemoryOrder = "Z  " ;
		QV_ADV_TEND:description = "tendency of qv adv" ;
		QV_ADV_TEND:units = "" ;
		QV_ADV_TEND:stagger = "" ;
		QV_ADV_TEND:_FillValue = -999.f ;
	float QV_RLX_TEND(Time, force_layers) ;
		QV_RLX_TEND:FieldType = 104 ;
		QV_RLX_TEND:MemoryOrder = "Z  " ;
		QV_RLX_TEND:description = "qv relaxation" ;
		QV_RLX_TEND:units = "" ;
		QV_RLX_TEND:stagger = "" ;
		QV_RLX_TEND:_FillValue = -999.f ;
        float INV_TAU_S(Time, force_layers) ;
                INV_TAU_S:FieldType = 104 ;
                INV_TAU_S:MemoryOrder = "Z  " ;
                INV_TAU_S:description = "inverse relaxation time for scalar" ;
                INV_TAU_S:units = "" ;
                INV_TAU_S:stagger = "" ;
                INV_TAU_S:_FillValue = -999.f ;
        float INV_TAU_M(Time, force_layers) ;
                INV_TAU_M:FieldType = 104 ;
                INV_TAU_M:MemoryOrder = "Z  " ;
                INV_TAU_M:description = "inverse relaxation time for momentum" ;
                INV_TAU_M:units = "" ;
                INV_TAU_M:stagger = "" ;
                INV_TAU_M:_FillValue = -999.f ;

// global attributes:
                :TITLE = "AUXILIARY FORCING FOR CRM" ;
}
